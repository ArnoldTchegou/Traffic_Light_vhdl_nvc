library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package constantes is
    constant Horloge : time := 1 ms; --paramétrable pour le testbench
end package constantes;
